oscillator_inst : oscillator PORT MAP (
		oscena	 => oscena_sig,
		osc	 => osc_sig
	);
